class sequence_item #(parameter width=8);
	rand logic [width-1:0]	in1;
	rand logic [width-1:0]	in0;
	     logic [width-1:0]	sum_out;
	     logic		carry_out;

	     function new();
	     endfunction 

endclass : sequence_item
